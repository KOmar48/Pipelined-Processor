`timescale 1ns / 1ps
/*
    AND module buh
*/
module AND (input AN0, AN1,
            output ANO);
            
assign ANO = AN0 & AN1;

endmodule
